magic
tech scmos
timestamp 1613667928
<< metal1 >>
rect -24 23 0 27
rect 992 23 1006 27
rect -24 -3 -20 23
rect 1002 -3 1006 23
rect -24 -7 1006 -3
use 5inv  5inv_0 5inv
timestamp 1613664914
transform 1 0 10 0 1 34
box -10 -34 22 35
use 5inv  5inv_1
timestamp 1613664914
transform 1 0 42 0 1 34
box -10 -34 22 35
use 5inv  5inv_2
timestamp 1613664914
transform 1 0 74 0 1 34
box -10 -34 22 35
use 5inv  5inv_3
timestamp 1613664914
transform 1 0 106 0 1 34
box -10 -34 22 35
use 5inv  5inv_4
timestamp 1613664914
transform 1 0 138 0 1 34
box -10 -34 22 35
use 5inv  5inv_5
timestamp 1613664914
transform 1 0 170 0 1 34
box -10 -34 22 35
use 5inv  5inv_6
timestamp 1613664914
transform 1 0 202 0 1 34
box -10 -34 22 35
use 5inv  5inv_7
timestamp 1613664914
transform 1 0 234 0 1 34
box -10 -34 22 35
use 5inv  5inv_8
timestamp 1613664914
transform 1 0 266 0 1 34
box -10 -34 22 35
use 5inv  5inv_9
timestamp 1613664914
transform 1 0 298 0 1 34
box -10 -34 22 35
use 5inv  5inv_10
timestamp 1613664914
transform 1 0 330 0 1 34
box -10 -34 22 35
use 5inv  5inv_11
timestamp 1613664914
transform 1 0 362 0 1 34
box -10 -34 22 35
use 5inv  5inv_12
timestamp 1613664914
transform 1 0 394 0 1 34
box -10 -34 22 35
use 5inv  5inv_13
timestamp 1613664914
transform 1 0 426 0 1 34
box -10 -34 22 35
use 5inv  5inv_14
timestamp 1613664914
transform 1 0 458 0 1 34
box -10 -34 22 35
use 5inv  5inv_15
timestamp 1613664914
transform 1 0 490 0 1 34
box -10 -34 22 35
use 5inv  5inv_16
timestamp 1613664914
transform 1 0 522 0 1 34
box -10 -34 22 35
use 5inv  5inv_17
timestamp 1613664914
transform 1 0 554 0 1 34
box -10 -34 22 35
use 5inv  5inv_18
timestamp 1613664914
transform 1 0 586 0 1 34
box -10 -34 22 35
use 5inv  5inv_19
timestamp 1613664914
transform 1 0 618 0 1 34
box -10 -34 22 35
use 5inv  5inv_20
timestamp 1613664914
transform 1 0 650 0 1 34
box -10 -34 22 35
use 5inv  5inv_21
timestamp 1613664914
transform 1 0 682 0 1 34
box -10 -34 22 35
use 5inv  5inv_22
timestamp 1613664914
transform 1 0 714 0 1 34
box -10 -34 22 35
use 5inv  5inv_23
timestamp 1613664914
transform 1 0 746 0 1 34
box -10 -34 22 35
use 5inv  5inv_24
timestamp 1613664914
transform 1 0 778 0 1 34
box -10 -34 22 35
use 5inv  5inv_25
timestamp 1613664914
transform 1 0 810 0 1 34
box -10 -34 22 35
use 5inv  5inv_26
timestamp 1613664914
transform 1 0 842 0 1 34
box -10 -34 22 35
use 5inv  5inv_27
timestamp 1613664914
transform 1 0 874 0 1 34
box -10 -34 22 35
use 5inv  5inv_28
timestamp 1613664914
transform 1 0 906 0 1 34
box -10 -34 22 35
use 5inv  5inv_29
timestamp 1613664914
transform 1 0 938 0 1 34
box -10 -34 22 35
use 5inv  5inv_30
timestamp 1613664914
transform 1 0 970 0 1 34
box -10 -34 22 35
<< end >>
